module test;
  initial begin
    $display("Hello from Verilog!");
    $finish;
  end
endmodule
